-- hi foo!

