dec_threshold_inst : dec_threshold PORT MAP (
		result	 => result_sig
	);
