library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use std.textio.all;
use work.cw_data_types.all;


package str21_data is

constant ATWD_SIZE_IN : integer := 64;
type simu_atwd_data_type is array (integer range 0 to atwd_size_in - 1) of word32;

constant SIMU_DATA : simu_atwd_data_type := 
(
B"00000000000000100000000000000011",
B"00000000000001010000000000000011",
B"00000000001110000000000000010110",
B"00000000001111010000000001001000",
B"00000000000110000000000000100111",
B"00000000000010010000000000010000",
B"00000000000001110000000000000111",
B"00000000000000110000000000000100",
B"00000000000001000000000000000011",
B"00000000000000110000000000000011",
B"00000000000000100000000000000010",
B"00000000000001000000000000000010",
B"00000000000001000000000000000011",
B"00000000000001000000000000000010",
B"00000000000011010000000000000111",
B"00000000000010100000000000001100",
B"00000000000011010000000000001000",
B"00000000000101100000000000010100",
B"00000000000010110000000000010000",
B"00000000000001100000000000000110",
B"00000000000001000000000000000011",
B"00000000000000110000000000000011",
B"00000000000001000000000000000011",
B"00000000000000010000000000000010",
B"00000000000000000000000000000010",
B"00000000000000110000000000000010",
B"00000000000000010000000000000001",
B"00000000000000100000000000000010",
B"00000000000000110000000000000011",
B"00000000000000110000000000000010",
B"00000000000000100000000000000010",
B"00000000000000100000000000000010",
B"00000000000000100000000000000010",
B"00000000000000110000000000000010",
B"00000000000000110000000000000010",
B"00000000000000110000000000000011",
B"00000000000000110000000000000010",
B"00000000000000100000000000000011",
B"00000000000000010000000000000001",
B"00000000000000100000000000000010",
B"00000000000000100000000000000010",
B"00000000000001000000000000000011",
B"00000000000000110000000000000100",
B"00000000000000110000000000000010",
B"00000000000000010000000000000011",
B"00000000000000100000000000000001",
B"00000000000000100000000000000001",
B"00000000000000110000000000000001",
B"00000000000001000000000000000010",
B"00000000000000110000000000000011",
B"00000000000000100000000000000010",
B"00000000000000110000000000000011",
B"00000000000000110000000000000011",
B"00000000000000110000000000000011",
B"00000000000000110000000000000011",
B"00000000000001010000000000000100",
B"00000000000000110000000000000100",
B"00000000000001000000000000000011",
B"00000000000000110000000000000011",
B"00000000000000010000000000000011",
B"00000000000000110000000000000010",
B"00000000000000110000000000000010",
B"00000000000000100000000000000001",
B"00000000000000110000000000000010"
);
end package;