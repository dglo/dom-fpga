-------------------------------------------------------------------------------
-- Title      : DOMAPP
-- Project    : IceCube DOM main board
-------------------------------------------------------------------------------
-- File       : compression.vhd
-- Author     : thorsten
-- Company    : LBNL
-- Created    : 
-- Last update: 2003-09-05
-- Platform   : Altera Excalibur
-- Standard   : VHDL'93
-------------------------------------------------------------------------------
-- Description: This module does the data compression on the ADC data
-------------------------------------------------------------------------------
-- Copyright (c) 2003 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version     Author    Description
-- 2003-09-05  V01-01-00   thorsten  
-------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.std_logic_arith.all;
USE IEEE.std_logic_unsigned.all;

USE WORK.icecube_data_types.all;
USE WORK.ctrl_data_types.all;

ENTITY compression IS
	GENERIC (
		FADC_WIDTH		: INTEGER := 10
		);
	PORT (
		CLK20		: IN STD_LOGIC;
		CLK40		: IN STD_LOGIC;
		RST			: IN STD_LOGIC;
		-- enable
		COMPR_ctrl	: IN COMPR_STRUCT;
		-- data input from data buffer
		data_avail_in	: IN STD_LOGIC;
		read_done_in	: OUT STD_LOGIC;
		HEADER_in		: IN HEADER_VECTOR;
		ATWD_addr_in	: OUT STD_LOGIC_VECTOR (7 downto 0);
		ATWD_data_in	: IN STD_LOGIC_VECTOR (31 downto 0);
		FADC_addr_in	: OUT STD_LOGIC_VECTOR (6 downto 0);
		FADC_data_in	: IN STD_LOGIC_VECTOR (31 downto 0);
		-- data output
		data_avail_out	: OUT STD_LOGIC;
		read_done_out	: IN STD_LOGIC;
		compr_avail_out	: OUT STD_LOGIC;
		compr_size		: OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
		compr_addr		: IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		compr_data		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
		HEADER_out		: OUT HEADER_VECTOR;
		ATWD_addr_out	: IN STD_LOGIC_VECTOR (7 downto 0);
		ATWD_data_out	: OUT STD_LOGIC_VECTOR (31 downto 0);
		FADC_addr_out	: IN STD_LOGIC_VECTOR (6 downto 0);
		FADC_data_out	: OUT STD_LOGIC_VECTOR (31 downto 0);
		-- test connector
		TC			: OUT STD_LOGIC_VECTOR(7 downto 0)
	);
END compression;


ARCHITECTURE arch_compression OF compression IS

BEGIN

	-- cpmression data
	--compr_avail_out <= '0';
	--compr_size		<= (OTHERS=>'0');
	compr_avail_out <= data_avail_in;
	compr_size		<= "111111011";
	PROCESS(CLK40)
	BEGIN
		IF CLK40'EVENT AND CLK40='1' THEN
			IF compr_addr=0 THEN
				compr_data <= x"deadbeef";
			ELSE
				compr_data (8 DOWNTO 0) <= compr_addr;
				compr_data (31 DOWNTO 9) <= (OTHERS=>'0');
				compr_data (24) <= '1';
			END IF;
		END IF;
	END PROCESS;
	
	--engineering data
	data_avail_out	<= data_avail_in;
	read_done_in	<= read_done_out;
	
	HEADER_out		<= HEADER_in;
	ATWD_addr_in	<= ATWD_addr_out;
	ATWD_data_out	<= ATWD_data_in;
	FADC_addr_in	<= FADC_addr_out;
	FADC_data_out	<= FADC_data_in;

END;
